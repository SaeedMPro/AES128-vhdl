library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Utilities is
    subtype BYTE is std_logic_vector(7 downto 0);
    type MATRIX is array (0 to 3,0 to 3) of BYTE;
    type stateOut is array (0 to 11) of MATRIX;
    type pipelineData is 
        record
            state: MATRIX;
            key: std_logic_vector(1407 downto 0);
            valid: std_logic;
        end record;
    type pipelineDataArray is array (0 to 10) of pipelineData;
    type roundKeyMatrix is array(0 to 10) of MATRIX;

    function plaintext_to_matrix(input_text: in std_logic_vector) return MATRIX;
    function matrix_to_plaintext(input_matrix: in MATRIX) return std_logic_vector;
    
    function two_mul_GF(input : BYTE) return BYTE;
    function mul_GF(input1 : BYTE; input2 : BYTE) return BYTE;
    
    function RotWord(word : std_logic_vector(31 downto 0)) return std_logic_vector;
    function SubWord(word : std_logic_vector(31 downto 0)) return std_logic_vector;

    constant mixColumn_matrix : MATRIX :=(
        (x"02", x"03", x"01", x"01"),
        (x"01", x"02", x"03", x"01"),
        (x"01", x"01", x"02", x"03"),
        (x"03", x"01", x"01", x"02")
    );
    constant inv_mixColumn_matrix : MATRIX := (
        (x"0E", x"0B", x"0D", x"09"),
        (x"09", x"0E", x"0B", x"0D"),
        (x"0D", x"09", x"0E", x"0B"),
        (x"0B", x"0D", x"09", x"0E")
    );

    type sbox_array is array (0 to 255) of std_logic_vector(7 downto 0);
    constant SBOX : sbox_array := (
        x"63", x"7C", x"77", x"7B", x"F2", x"6B", x"6F", x"C5",
        x"30", x"01", x"67", x"2B", x"FE", x"D7", x"AB", x"76",
        x"CA", x"82", x"C9", x"7D", x"FA", x"59", x"47", x"F0",
        x"AD", x"D4", x"A2", x"AF", x"9C", x"A4", x"72", x"C0",
        x"B7", x"FD", x"93", x"26", x"36", x"3F", x"F7", x"CC",
        x"34", x"A5", x"E5", x"F1", x"71", x"D8", x"31", x"15",
        x"04", x"C7", x"23", x"C3", x"18", x"96", x"05", x"9A",
        x"07", x"12", x"80", x"E2", x"EB", x"27", x"B2", x"75",
        x"09", x"83", x"2C", x"1A", x"1B", x"6E", x"5A", x"A0",
        x"52", x"3B", x"D6", x"B3", x"29", x"E3", x"2F", x"84",
        x"53", x"D1", x"00", x"ED", x"20", x"FC", x"B1", x"5B",
        x"6A", x"CB", x"BE", x"39", x"4A", x"4C", x"58", x"CF",
        x"D0", x"EF", x"AA", x"FB", x"43", x"4D", x"33", x"85",
        x"45", x"F9", x"02", x"7F", x"50", x"3C", x"9F", x"A8",
        x"51", x"A3", x"40", x"8F", x"92", x"9D", x"38", x"F5",
        x"BC", x"B6", x"DA", x"21", x"10", x"FF", x"F3", x"D2",
        x"CD", x"0C", x"13", x"EC", x"5F", x"97", x"44", x"17",
        x"C4", x"A7", x"7E", x"3D", x"64", x"5D", x"19", x"73",
        x"60", x"81", x"4F", x"DC", x"22", x"2A", x"90", x"88",
        x"46", x"EE", x"B8", x"14", x"DE", x"5E", x"0B", x"DB",
        x"E0", x"32", x"3A", x"0A", x"49", x"06", x"24", x"5C",
        x"C2", x"D3", x"AC", x"62", x"91", x"95", x"E4", x"79",
        x"E7", x"C8", x"37", x"6D", x"8D", x"D5", x"4E", x"A9",
        x"6C", x"56", x"F4", x"EA", x"65", x"7A", x"AE", x"08",
        x"BA", x"78", x"25", x"2E", x"1C", x"A6", x"B4", x"C6",
        x"E8", x"DD", x"74", x"1F", x"4B", x"BD", x"8B", x"8A",
        x"70", x"3E", x"B5", x"66", x"48", x"03", x"F6", x"0E",
        x"61", x"35", x"57", x"B9", x"86", x"C1", x"1D", x"9E",
        x"E1", x"F8", x"98", x"11", x"69", x"D9", x"8E", x"94",
        x"9B", x"1E", x"87", x"E9", x"CE", x"55", x"28", x"DF",
        x"8C", x"A1", x"89", x"0D", x"BF", x"E6", x"42", x"68",
        x"41", x"99", x"2D", x"0F", x"B0", x"54", x"BB", x"16"
    );
    constant INV_SBOX : sbox_array := (
        x"52", x"09", x"6A", x"D5", x"30", x"36", x"A5", x"38",
        x"BF", x"40", x"A3", x"9E", x"81", x"F3", x"D7", x"FB",
        x"7C", x"E3", x"39", x"82", x"9B", x"2F", x"FF", x"87",
        x"34", x"8E", x"43", x"44", x"C4", x"DE", x"E9", x"CB",
        x"54", x"7B", x"94", x"32", x"A6", x"C2", x"23", x"3D",
        x"EE", x"4C", x"95", x"0B", x"42", x"FA", x"C3", x"4E",
        x"08", x"2E", x"A1", x"66", x"28", x"D9", x"24", x"B2",
        x"76", x"5B", x"A2", x"49", x"6D", x"8B", x"D1", x"25",
        x"72", x"F8", x"F6", x"64", x"86", x"68", x"98", x"16",
        x"D4", x"A4", x"5C", x"CC", x"5D", x"65", x"B6", x"92",
        x"6C", x"70", x"48", x"50", x"FD", x"ED", x"B9", x"DA",
        x"5E", x"15", x"46", x"57", x"A7", x"8D", x"9D", x"84",
        x"90", x"D8", x"AB", x"00", x"8C", x"BC", x"D3", x"0A",
        x"F7", x"E4", x"58", x"05", x"B8", x"B3", x"45", x"06",
        x"D0", x"2C", x"1E", x"8F", x"CA", x"3F", x"0F", x"02",
        x"C1", x"AF", x"BD", x"03", x"01", x"13", x"8A", x"6B",
        x"3A", x"91", x"11", x"41", x"4F", x"67", x"DC", x"EA",
        x"97", x"F2", x"CF", x"CE", x"F0", x"B4", x"E6", x"73",
        x"96", x"AC", x"74", x"22", x"E7", x"AD", x"35", x"85",
        x"E2", x"F9", x"37", x"E8", x"1C", x"75", x"DF", x"6E",
        x"47", x"F1", x"1A", x"71", x"1D", x"29", x"C5", x"89",
        x"6F", x"B7", x"62", x"0E", x"AA", x"18", x"BE", x"1B",
        x"FC", x"56", x"3E", x"4B", x"C6", x"D2", x"79", x"20",
        x"9A", x"DB", x"C0", x"FE", x"78", x"CD", x"5A", x"F4",
        x"1F", x"DD", x"A8", x"33", x"88", x"07", x"C7", x"31",
        x"B1", x"12", x"10", x"59", x"27", x"80", x"EC", x"5F",
        x"60", x"51", x"7F", x"A9", x"19", x"B5", x"4A", x"0D",
        x"2D", x"E5", x"7A", x"9F", x"93", x"C9", x"9C", x"EF",
        x"A0", x"E0", x"3B", x"4D", x"AE", x"2A", x"F5", x"B0",
        x"C8", x"EB", x"BB", x"3C", x"83", x"53", x"99", x"61",
        x"17", x"2B", x"04", x"7E", x"BA", x"77", x"D6", x"26",
        x"E1", x"69", x"14", x"63", x"55", x"21", x"0C", x"7D"
    );

    type rcon_array is array(0 to 10) of std_logic_vector(31 downto 0);
    constant RCON : rcon_array := (
        x"01000000", x"02000000", x"04000000", x"08000000", x"10000000",
        x"20000000", x"40000000", x"80000000", x"1B000000", x"36000000", x"00000000"
    );
        
 end Utilities;

package body Utilities is

    function plaintext_to_matrix(input_text: in std_logic_vector) return MATRIX is
        variable output_matrix: MATRIX;
    begin
        for j in 3 downto 0 loop 
                for i in 3 downto 0 loop
                    output_matrix(i,j) := input_text(input_text'high-(j*32 + i*8) downto (input_text'high-(j*32 + i*8))-7);
                end loop;
        end loop;
        return output_matrix;
    end function;

    function matrix_to_plaintext(input_matrix: in MATRIX) return std_logic_vector is
        variable output_text: std_logic_vector(127 downto 0);
    begin
        for j in 3 downto 0 loop 
			for i in 3 downto 0 loop
				output_text(127-(j*32 + i*8) downto (127-(j*32 + i*8))-7) := input_matrix(i,j);
			end loop;
        end loop;
        return output_text;
    end function;

    function RotWord(word : std_logic_vector(31 downto 0)) return std_logic_vector is
        variable w : std_logic_vector(31 downto 0);
    begin
        w := word(23 downto 0) & word(31 downto 24);
        return w;
    end function;

    function SubWord(word : std_logic_vector(31 downto 0)) return std_logic_vector is
        variable w : std_logic_vector(31 downto 0);
    begin
        for i in 0 to 3 loop
                w(8*(3-i)+7 downto 8*(3-i)) := SBOX(to_integer(unsigned(word(8*(3-i)+7 downto 8*(3-i)))));
        end loop;
        return w;
    end function;

    function two_mul_GF(input : BYTE) return BYTE is
        variable shifted : BYTE := (others => '0');
        variable result  : BYTE := (others => '0');
    begin
        shifted := input(6 downto 0) & '0';
        if input(7) = '1' then
            result := shifted xor x"1B";
        else
            result := shifted;
        end if;
        return result;
    end function;

	function mul_GF(input1 : BYTE; input2 : BYTE) return BYTE is
        variable t1, t2, t3, res : BYTE := (others => '0');
	begin
        case input2 is
            when x"01" =>
                res := input1;
            when x"02" =>
                res := two_mul_GF(input1);
            when x"03" =>
                res := std_logic_vector(unsigned(two_mul_GF(input1)) xor unsigned(input1));
            when x"09" =>
                t1 := two_mul_GF(input1);
                t2 := two_mul_GF(t1);
                t3 := two_mul_GF(t2);
                res := std_logic_vector(unsigned(t3) xor unsigned(input1));
            when x"0B" =>
                t1 := two_mul_GF(input1);      
                t2 := two_mul_GF(t1);     
                t3 := two_mul_GF(t2);     
                res := std_logic_vector(unsigned(t3) xor unsigned(t1) xor unsigned(input1));
            when x"0D" =>
                t1 := two_mul_GF(input1);      
                t2 := two_mul_GF(t1);     
                t3 := two_mul_GF(t2);     
                res := std_logic_vector(unsigned(t3) xor unsigned(t2) xor unsigned(input1));
            when x"0E" =>
                t1 := two_mul_GF(input1);      
                t2 := two_mul_GF(t1);     
                t3 := two_mul_GF(t2);     
                res := std_logic_vector(unsigned(t3) xor unsigned(t2) xor unsigned(t1));
            when others =>
                res := (others => '0');
        end case;
        return res;
	end function;

end Utilities;
