
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Utilities is

 SUBTYPE WORD_8BIT IS STD_LOGIC_VECTOR(7 DOWNTO 0);
 TYPE MATRIX IS ARRAY (0 TO 3,0 TO 3) OF WORD_8BIT;

end Utilities;

package body Utilities is
 
end Utilities;
