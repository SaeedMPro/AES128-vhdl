library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity shiftrows is
end shiftrows;

architecture Behavioral of shiftrows is
begin

end Behavioral;
