library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity sbox is
    Port (

        );
end sbox;

architecture Behavioral of sbox is
begin

end Behavioral;
