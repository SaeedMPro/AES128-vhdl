library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity mixcolumns is
    Port (

        );
end mixcolumns;

architecture Behavioral of mixcolumns is
begin

end Behavioral;
