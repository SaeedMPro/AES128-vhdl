library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity subbytes is
    Port (

        );
end subbytes;

architecture Behavioral of subbytes is
begin

end Behavioral;
