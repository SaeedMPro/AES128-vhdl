library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity addroundkey is
    Port (
        
        );
end addroundkey;

architecture Behavioral of addroundkey is
begin

end Behavioral;
